module add4(
    input [31:0] pcOut,
    output [31:0] add4Out
);
    
    assign add4Out = pcOut + 4;

endmodule
