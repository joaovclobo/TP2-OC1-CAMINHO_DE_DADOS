module add4(
    input [31:0] pcIn,
    output [31:0] add4
);
    
    assign add4 = pcIn + 4;

endmodule
